library verilog;
use verilog.vl_types.all;
entity T_flipflop_vlg_vec_tst is
end T_flipflop_vlg_vec_tst;
