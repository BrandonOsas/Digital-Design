library verilog;
use verilog.vl_types.all;
entity Gray_code4_vlg_vec_tst is
end Gray_code4_vlg_vec_tst;
