library verilog;
use verilog.vl_types.all;
entity LAb1_vlg_vec_tst is
end LAb1_vlg_vec_tst;
