library verilog;
use verilog.vl_types.all;
entity Taillight_vlg_vec_tst is
end Taillight_vlg_vec_tst;
