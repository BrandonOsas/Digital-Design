library verilog;
use verilog.vl_types.all;
entity counter16_vlg_vec_tst is
end counter16_vlg_vec_tst;
